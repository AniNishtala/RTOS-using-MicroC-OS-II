// unsaved.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module unsaved (
		input  wire        clk_clk,         //        clk.clk
		output wire [6:0]  hex0_export,     //       hex0.export
		output wire [6:0]  hex1_export,     //       hex1.export
		output wire [6:0]  hex2_export,     //       hex2.export
		output wire [6:0]  hex3_export,     //       hex3.export
		output wire [6:0]  hex4_export,     //       hex4.export
		output wire [6:0]  hex5_export,     //       hex5.export
		output wire [6:0]  hex6_export,     //       hex6.export
		output wire [6:0]  hex7_export,     //       hex7.export
		output wire [31:0] jp5_export,      //        jp5.export
		input  wire [2:0]  key_export,      //        key.export
		inout  wire [7:0]  lcd_module_DATA, // lcd_module.DATA
		output wire        lcd_module_ON,   //           .ON
		output wire        lcd_module_BLON, //           .BLON
		output wire        lcd_module_EN,   //           .EN
		output wire        lcd_module_RS,   //           .RS
		output wire        lcd_module_RW,   //           .RW
		output wire [7:0]  ledg_export,     //       ledg.export
		output wire [17:0] ledr_export,     //       ledr.export
		input  wire        reset_reset,     //      reset.reset
		output wire [11:0] sdram_addr,      //      sdram.addr
		output wire [1:0]  sdram_ba,        //           .ba
		output wire        sdram_cas_n,     //           .cas_n
		output wire        sdram_cke,       //           .cke
		output wire        sdram_cs_n,      //           .cs_n
		inout  wire [31:0] sdram_dq,        //           .dq
		output wire [3:0]  sdram_dqm,       //           .dqm
		output wire        sdram_ras_n,     //           .ras_n
		output wire        sdram_we_n,      //           .we_n
		output wire        sdram_clk_clk,   //  sdram_clk.clk
		inout  wire [15:0] sram_DQ,         //       sram.DQ
		output wire [19:0] sram_ADDR,       //           .ADDR
		output wire        sram_LB_N,       //           .LB_N
		output wire        sram_UB_N,       //           .UB_N
		output wire        sram_CE_N,       //           .CE_N
		output wire        sram_OE_N,       //           .OE_N
		output wire        sram_WE_N,       //           .WE_N
		input  wire [17:0] switches_export  //   switches.export
	);

	wire         clocks_sys_clk_clk;                                           // clocks:sys_clk_clk -> [GPIO:clk, HEX0:clk, HEX1:clk, HEX2:clk, HEX3:clk, HEX4:clk, HEX5:clk, HEX6:clk, HEX7:clk, HIGH_TIMER:clk, KEY:clk, LCD_DATA:clk, LEDG:clk, LEDR:clk, SW:clk, SYSTEM_TIMER:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:clocks_sys_clk_clk, nios2_qsys_0:clk, on_chip_memory:clk, rst_controller:clk, sdram:clk, sram:clk, sysid_qsys_0:clock]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> [GPIO:reset_n, LCD_DATA:reset, mm_interconnect_0:LCD_DATA_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [25:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [25:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_lcd_data_avalon_lcd_slave_chipselect;       // mm_interconnect_0:LCD_DATA_avalon_lcd_slave_chipselect -> LCD_DATA:chipselect
	wire   [7:0] mm_interconnect_0_lcd_data_avalon_lcd_slave_readdata;         // LCD_DATA:readdata -> mm_interconnect_0:LCD_DATA_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_lcd_data_avalon_lcd_slave_waitrequest;      // LCD_DATA:waitrequest -> mm_interconnect_0:LCD_DATA_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_lcd_data_avalon_lcd_slave_address;          // mm_interconnect_0:LCD_DATA_avalon_lcd_slave_address -> LCD_DATA:address
	wire         mm_interconnect_0_lcd_data_avalon_lcd_slave_read;             // mm_interconnect_0:LCD_DATA_avalon_lcd_slave_read -> LCD_DATA:read
	wire         mm_interconnect_0_lcd_data_avalon_lcd_slave_write;            // mm_interconnect_0:LCD_DATA_avalon_lcd_slave_write -> LCD_DATA:write
	wire   [7:0] mm_interconnect_0_lcd_data_avalon_lcd_slave_writedata;        // mm_interconnect_0:LCD_DATA_avalon_lcd_slave_writedata -> LCD_DATA:writedata
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;            // sram:readdata -> mm_interconnect_0:sram_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;             // mm_interconnect_0:sram_avalon_sram_slave_address -> sram:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                // mm_interconnect_0:sram_avalon_sram_slave_read -> sram:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;          // mm_interconnect_0:sram_avalon_sram_slave_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;       // sram:readdatavalid -> mm_interconnect_0:sram_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;               // mm_interconnect_0:sram_avalon_sram_slave_write -> sram:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;           // mm_interconnect_0:sram_avalon_sram_slave_writedata -> sram:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;        // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;         // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_on_chip_memory_s1_chipselect;               // mm_interconnect_0:on_chip_memory_s1_chipselect -> on_chip_memory:chipselect
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_readdata;                 // on_chip_memory:readdata -> mm_interconnect_0:on_chip_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_on_chip_memory_s1_address;                  // mm_interconnect_0:on_chip_memory_s1_address -> on_chip_memory:address
	wire   [3:0] mm_interconnect_0_on_chip_memory_s1_byteenable;               // mm_interconnect_0:on_chip_memory_s1_byteenable -> on_chip_memory:byteenable
	wire         mm_interconnect_0_on_chip_memory_s1_write;                    // mm_interconnect_0:on_chip_memory_s1_write -> on_chip_memory:write
	wire  [31:0] mm_interconnect_0_on_chip_memory_s1_writedata;                // mm_interconnect_0:on_chip_memory_s1_writedata -> on_chip_memory:writedata
	wire         mm_interconnect_0_on_chip_memory_s1_clken;                    // mm_interconnect_0:on_chip_memory_s1_clken -> on_chip_memory:clken
	wire         mm_interconnect_0_sw_s1_chipselect;                           // mm_interconnect_0:SW_s1_chipselect -> SW:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                             // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                              // mm_interconnect_0:SW_s1_address -> SW:address
	wire         mm_interconnect_0_sw_s1_write;                                // mm_interconnect_0:SW_s1_write -> SW:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                            // mm_interconnect_0:SW_s1_writedata -> SW:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                         // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                           // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                            // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                              // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                          // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_ledg_s1_chipselect;                         // mm_interconnect_0:LEDG_s1_chipselect -> LEDG:chipselect
	wire  [31:0] mm_interconnect_0_ledg_s1_readdata;                           // LEDG:readdata -> mm_interconnect_0:LEDG_s1_readdata
	wire   [1:0] mm_interconnect_0_ledg_s1_address;                            // mm_interconnect_0:LEDG_s1_address -> LEDG:address
	wire         mm_interconnect_0_ledg_s1_write;                              // mm_interconnect_0:LEDG_s1_write -> LEDG:write_n
	wire  [31:0] mm_interconnect_0_ledg_s1_writedata;                          // mm_interconnect_0:LEDG_s1_writedata -> LEDG:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                          // mm_interconnect_0:KEY_s1_chipselect -> KEY:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                            // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                             // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_key_s1_write;                               // mm_interconnect_0:KEY_s1_write -> KEY:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                           // mm_interconnect_0:KEY_s1_writedata -> KEY:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                         // mm_interconnect_0:HEX0_s1_chipselect -> HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                           // HEX0:readdata -> mm_interconnect_0:HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                            // mm_interconnect_0:HEX0_s1_address -> HEX0:address
	wire         mm_interconnect_0_hex0_s1_write;                              // mm_interconnect_0:HEX0_s1_write -> HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                          // mm_interconnect_0:HEX0_s1_writedata -> HEX0:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                         // mm_interconnect_0:HEX1_s1_chipselect -> HEX1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                           // HEX1:readdata -> mm_interconnect_0:HEX1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                            // mm_interconnect_0:HEX1_s1_address -> HEX1:address
	wire         mm_interconnect_0_hex1_s1_write;                              // mm_interconnect_0:HEX1_s1_write -> HEX1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                          // mm_interconnect_0:HEX1_s1_writedata -> HEX1:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                         // mm_interconnect_0:HEX2_s1_chipselect -> HEX2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                           // HEX2:readdata -> mm_interconnect_0:HEX2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                            // mm_interconnect_0:HEX2_s1_address -> HEX2:address
	wire         mm_interconnect_0_hex2_s1_write;                              // mm_interconnect_0:HEX2_s1_write -> HEX2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                          // mm_interconnect_0:HEX2_s1_writedata -> HEX2:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                         // mm_interconnect_0:HEX3_s1_chipselect -> HEX3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                           // HEX3:readdata -> mm_interconnect_0:HEX3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                            // mm_interconnect_0:HEX3_s1_address -> HEX3:address
	wire         mm_interconnect_0_hex3_s1_write;                              // mm_interconnect_0:HEX3_s1_write -> HEX3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                          // mm_interconnect_0:HEX3_s1_writedata -> HEX3:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                         // mm_interconnect_0:HEX4_s1_chipselect -> HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                           // HEX4:readdata -> mm_interconnect_0:HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                            // mm_interconnect_0:HEX4_s1_address -> HEX4:address
	wire         mm_interconnect_0_hex4_s1_write;                              // mm_interconnect_0:HEX4_s1_write -> HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                          // mm_interconnect_0:HEX4_s1_writedata -> HEX4:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                         // mm_interconnect_0:HEX5_s1_chipselect -> HEX5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                           // HEX5:readdata -> mm_interconnect_0:HEX5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                            // mm_interconnect_0:HEX5_s1_address -> HEX5:address
	wire         mm_interconnect_0_hex5_s1_write;                              // mm_interconnect_0:HEX5_s1_write -> HEX5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                          // mm_interconnect_0:HEX5_s1_writedata -> HEX5:writedata
	wire         mm_interconnect_0_hex6_s1_chipselect;                         // mm_interconnect_0:HEX6_s1_chipselect -> HEX6:chipselect
	wire  [31:0] mm_interconnect_0_hex6_s1_readdata;                           // HEX6:readdata -> mm_interconnect_0:HEX6_s1_readdata
	wire   [1:0] mm_interconnect_0_hex6_s1_address;                            // mm_interconnect_0:HEX6_s1_address -> HEX6:address
	wire         mm_interconnect_0_hex6_s1_write;                              // mm_interconnect_0:HEX6_s1_write -> HEX6:write_n
	wire  [31:0] mm_interconnect_0_hex6_s1_writedata;                          // mm_interconnect_0:HEX6_s1_writedata -> HEX6:writedata
	wire         mm_interconnect_0_hex7_s1_chipselect;                         // mm_interconnect_0:HEX7_s1_chipselect -> HEX7:chipselect
	wire  [31:0] mm_interconnect_0_hex7_s1_readdata;                           // HEX7:readdata -> mm_interconnect_0:HEX7_s1_readdata
	wire   [1:0] mm_interconnect_0_hex7_s1_address;                            // mm_interconnect_0:HEX7_s1_address -> HEX7:address
	wire         mm_interconnect_0_hex7_s1_write;                              // mm_interconnect_0:HEX7_s1_write -> HEX7:write_n
	wire  [31:0] mm_interconnect_0_hex7_s1_writedata;                          // mm_interconnect_0:HEX7_s1_writedata -> HEX7:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_system_timer_s1_chipselect;                 // mm_interconnect_0:SYSTEM_TIMER_s1_chipselect -> SYSTEM_TIMER:chipselect
	wire  [15:0] mm_interconnect_0_system_timer_s1_readdata;                   // SYSTEM_TIMER:readdata -> mm_interconnect_0:SYSTEM_TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_system_timer_s1_address;                    // mm_interconnect_0:SYSTEM_TIMER_s1_address -> SYSTEM_TIMER:address
	wire         mm_interconnect_0_system_timer_s1_write;                      // mm_interconnect_0:SYSTEM_TIMER_s1_write -> SYSTEM_TIMER:write_n
	wire  [15:0] mm_interconnect_0_system_timer_s1_writedata;                  // mm_interconnect_0:SYSTEM_TIMER_s1_writedata -> SYSTEM_TIMER:writedata
	wire         mm_interconnect_0_high_timer_s1_chipselect;                   // mm_interconnect_0:HIGH_TIMER_s1_chipselect -> HIGH_TIMER:chipselect
	wire  [15:0] mm_interconnect_0_high_timer_s1_readdata;                     // HIGH_TIMER:readdata -> mm_interconnect_0:HIGH_TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_high_timer_s1_address;                      // mm_interconnect_0:HIGH_TIMER_s1_address -> HIGH_TIMER:address
	wire         mm_interconnect_0_high_timer_s1_write;                        // mm_interconnect_0:HIGH_TIMER_s1_write -> HIGH_TIMER:write_n
	wire  [15:0] mm_interconnect_0_high_timer_s1_writedata;                    // mm_interconnect_0:HIGH_TIMER_s1_writedata -> HIGH_TIMER:writedata
	wire         mm_interconnect_0_gpio_s1_chipselect;                         // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;                           // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;                            // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;                              // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;                          // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         irq_mapper_receiver0_irq;                                     // KEY:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // SYSTEM_TIMER:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                     // HIGH_TIMER:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                     // SW:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [HEX0:reset_n, HEX1:reset_n, HEX2:reset_n, HEX3:reset_n, HEX4:reset_n, HEX5:reset_n, HEX6:reset_n, HEX7:reset_n, HIGH_TIMER:reset_n, KEY:reset_n, LEDG:reset_n, LEDR:reset_n, SW:reset_n, SYSTEM_TIMER:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, on_chip_memory:reset, rst_translator:in_reset, sdram:reset_n, sram:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, on_chip_memory:reset_req, rst_translator:reset_req_in]
	wire         clocks_reset_source_reset;                                    // clocks:reset_source_reset -> rst_controller:reset_in1

	unsaved_GPIO gpio (
		.clk        (clocks_sys_clk_clk),                          //                 clk.clk
		.reset_n    (~nios2_qsys_0_jtag_debug_module_reset_reset), //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),           //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),            //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),         //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect),        //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),          //                    .readdata
		.out_port   (jp5_export)                                   // external_connection.export
	);

	unsaved_HEX0 hex0 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                           // external_connection.export
	);

	unsaved_HEX0 hex1 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                           // external_connection.export
	);

	unsaved_HEX0 hex2 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                           // external_connection.export
	);

	unsaved_HEX0 hex3 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                           // external_connection.export
	);

	unsaved_HEX0 hex4 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                           // external_connection.export
	);

	unsaved_HEX0 hex5 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                           // external_connection.export
	);

	unsaved_HEX0 hex6 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex6_s1_readdata),   //                    .readdata
		.out_port   (hex6_export)                           // external_connection.export
	);

	unsaved_HEX0 hex7 (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex7_s1_readdata),   //                    .readdata
		.out_port   (hex7_export)                           // external_connection.export
	);

	unsaved_HIGH_TIMER high_timer (
		.clk        (clocks_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            // reset.reset_n
		.address    (mm_interconnect_0_high_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_high_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_high_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_high_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_high_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                    //   irq.irq
	);

	unsaved_KEY key (
		.clk        (clocks_sys_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_export),                          // external_connection.export
		.irq        (irq_mapper_receiver0_irq)             //                 irq.irq
	);

	unsaved_LCD_DATA lcd_data (
		.clk         (clocks_sys_clk_clk),                                      //                clk.clk
		.reset       (nios2_qsys_0_jtag_debug_module_reset_reset),              //              reset.reset
		.address     (mm_interconnect_0_lcd_data_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_lcd_data_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_lcd_data_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_lcd_data_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_lcd_data_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_lcd_data_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_lcd_data_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_module_DATA),                                         // external_interface.export
		.LCD_ON      (lcd_module_ON),                                           //                   .export
		.LCD_BLON    (lcd_module_BLON),                                         //                   .export
		.LCD_EN      (lcd_module_EN),                                           //                   .export
		.LCD_RS      (lcd_module_RS),                                           //                   .export
		.LCD_RW      (lcd_module_RW)                                            //                   .export
	);

	unsaved_LEDG ledg (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledg_s1_readdata),   //                    .readdata
		.out_port   (ledg_export)                           // external_connection.export
	);

	unsaved_LEDR ledr (
		.clk        (clocks_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	unsaved_SW sw (
		.clk        (clocks_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (switches_export),                    // external_connection.export
		.irq        (irq_mapper_receiver4_irq)            //                 irq.irq
	);

	unsaved_SYSTEM_TIMER system_timer (
		.clk        (clocks_sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_system_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_system_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_system_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_system_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_system_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                      //   irq.irq
	);

	unsaved_clocks clocks (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (reset_reset),               //    ref_reset.reset
		.sys_clk_clk        (clocks_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),             //    sdram_clk.clk
		.reset_source_reset (clocks_reset_source_reset)  // reset_source.reset
	);

	unsaved_jtag_uart_0 jtag_uart_0 (
		.clk            (clocks_sys_clk_clk),                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	unsaved_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clocks_sys_clk_clk),                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	unsaved_on_chip_memory on_chip_memory (
		.clk        (clocks_sys_clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_on_chip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_on_chip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_on_chip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_on_chip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_on_chip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_on_chip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_on_chip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	unsaved_sdram sdram (
		.clk            (clocks_sys_clk_clk),                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	unsaved_sram sram (
		.clk           (clocks_sys_clk_clk),                                     //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                              //                   .export
		.SRAM_LB_N     (sram_LB_N),                                              //                   .export
		.SRAM_UB_N     (sram_UB_N),                                              //                   .export
		.SRAM_CE_N     (sram_CE_N),                                              //                   .export
		.SRAM_OE_N     (sram_OE_N),                                              //                   .export
		.SRAM_WE_N     (sram_WE_N),                                              //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	unsaved_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clocks_sys_clk_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	unsaved_mm_interconnect_0 mm_interconnect_0 (
		.clocks_sys_clk_clk                               (clocks_sys_clk_clk),                                           //                             clocks_sys_clk.clk
		.LCD_DATA_reset_reset_bridge_in_reset_reset       (nios2_qsys_0_jtag_debug_module_reset_reset),                   //       LCD_DATA_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_readdatavalid           (nios2_qsys_0_data_master_readdatavalid),                       //                                           .readdatavalid
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.nios2_qsys_0_instruction_master_readdatavalid    (nios2_qsys_0_instruction_master_readdatavalid),                //                                           .readdatavalid
		.GPIO_s1_address                                  (mm_interconnect_0_gpio_s1_address),                            //                                    GPIO_s1.address
		.GPIO_s1_write                                    (mm_interconnect_0_gpio_s1_write),                              //                                           .write
		.GPIO_s1_readdata                                 (mm_interconnect_0_gpio_s1_readdata),                           //                                           .readdata
		.GPIO_s1_writedata                                (mm_interconnect_0_gpio_s1_writedata),                          //                                           .writedata
		.GPIO_s1_chipselect                               (mm_interconnect_0_gpio_s1_chipselect),                         //                                           .chipselect
		.HEX0_s1_address                                  (mm_interconnect_0_hex0_s1_address),                            //                                    HEX0_s1.address
		.HEX0_s1_write                                    (mm_interconnect_0_hex0_s1_write),                              //                                           .write
		.HEX0_s1_readdata                                 (mm_interconnect_0_hex0_s1_readdata),                           //                                           .readdata
		.HEX0_s1_writedata                                (mm_interconnect_0_hex0_s1_writedata),                          //                                           .writedata
		.HEX0_s1_chipselect                               (mm_interconnect_0_hex0_s1_chipselect),                         //                                           .chipselect
		.HEX1_s1_address                                  (mm_interconnect_0_hex1_s1_address),                            //                                    HEX1_s1.address
		.HEX1_s1_write                                    (mm_interconnect_0_hex1_s1_write),                              //                                           .write
		.HEX1_s1_readdata                                 (mm_interconnect_0_hex1_s1_readdata),                           //                                           .readdata
		.HEX1_s1_writedata                                (mm_interconnect_0_hex1_s1_writedata),                          //                                           .writedata
		.HEX1_s1_chipselect                               (mm_interconnect_0_hex1_s1_chipselect),                         //                                           .chipselect
		.HEX2_s1_address                                  (mm_interconnect_0_hex2_s1_address),                            //                                    HEX2_s1.address
		.HEX2_s1_write                                    (mm_interconnect_0_hex2_s1_write),                              //                                           .write
		.HEX2_s1_readdata                                 (mm_interconnect_0_hex2_s1_readdata),                           //                                           .readdata
		.HEX2_s1_writedata                                (mm_interconnect_0_hex2_s1_writedata),                          //                                           .writedata
		.HEX2_s1_chipselect                               (mm_interconnect_0_hex2_s1_chipselect),                         //                                           .chipselect
		.HEX3_s1_address                                  (mm_interconnect_0_hex3_s1_address),                            //                                    HEX3_s1.address
		.HEX3_s1_write                                    (mm_interconnect_0_hex3_s1_write),                              //                                           .write
		.HEX3_s1_readdata                                 (mm_interconnect_0_hex3_s1_readdata),                           //                                           .readdata
		.HEX3_s1_writedata                                (mm_interconnect_0_hex3_s1_writedata),                          //                                           .writedata
		.HEX3_s1_chipselect                               (mm_interconnect_0_hex3_s1_chipselect),                         //                                           .chipselect
		.HEX4_s1_address                                  (mm_interconnect_0_hex4_s1_address),                            //                                    HEX4_s1.address
		.HEX4_s1_write                                    (mm_interconnect_0_hex4_s1_write),                              //                                           .write
		.HEX4_s1_readdata                                 (mm_interconnect_0_hex4_s1_readdata),                           //                                           .readdata
		.HEX4_s1_writedata                                (mm_interconnect_0_hex4_s1_writedata),                          //                                           .writedata
		.HEX4_s1_chipselect                               (mm_interconnect_0_hex4_s1_chipselect),                         //                                           .chipselect
		.HEX5_s1_address                                  (mm_interconnect_0_hex5_s1_address),                            //                                    HEX5_s1.address
		.HEX5_s1_write                                    (mm_interconnect_0_hex5_s1_write),                              //                                           .write
		.HEX5_s1_readdata                                 (mm_interconnect_0_hex5_s1_readdata),                           //                                           .readdata
		.HEX5_s1_writedata                                (mm_interconnect_0_hex5_s1_writedata),                          //                                           .writedata
		.HEX5_s1_chipselect                               (mm_interconnect_0_hex5_s1_chipselect),                         //                                           .chipselect
		.HEX6_s1_address                                  (mm_interconnect_0_hex6_s1_address),                            //                                    HEX6_s1.address
		.HEX6_s1_write                                    (mm_interconnect_0_hex6_s1_write),                              //                                           .write
		.HEX6_s1_readdata                                 (mm_interconnect_0_hex6_s1_readdata),                           //                                           .readdata
		.HEX6_s1_writedata                                (mm_interconnect_0_hex6_s1_writedata),                          //                                           .writedata
		.HEX6_s1_chipselect                               (mm_interconnect_0_hex6_s1_chipselect),                         //                                           .chipselect
		.HEX7_s1_address                                  (mm_interconnect_0_hex7_s1_address),                            //                                    HEX7_s1.address
		.HEX7_s1_write                                    (mm_interconnect_0_hex7_s1_write),                              //                                           .write
		.HEX7_s1_readdata                                 (mm_interconnect_0_hex7_s1_readdata),                           //                                           .readdata
		.HEX7_s1_writedata                                (mm_interconnect_0_hex7_s1_writedata),                          //                                           .writedata
		.HEX7_s1_chipselect                               (mm_interconnect_0_hex7_s1_chipselect),                         //                                           .chipselect
		.HIGH_TIMER_s1_address                            (mm_interconnect_0_high_timer_s1_address),                      //                              HIGH_TIMER_s1.address
		.HIGH_TIMER_s1_write                              (mm_interconnect_0_high_timer_s1_write),                        //                                           .write
		.HIGH_TIMER_s1_readdata                           (mm_interconnect_0_high_timer_s1_readdata),                     //                                           .readdata
		.HIGH_TIMER_s1_writedata                          (mm_interconnect_0_high_timer_s1_writedata),                    //                                           .writedata
		.HIGH_TIMER_s1_chipselect                         (mm_interconnect_0_high_timer_s1_chipselect),                   //                                           .chipselect
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.KEY_s1_address                                   (mm_interconnect_0_key_s1_address),                             //                                     KEY_s1.address
		.KEY_s1_write                                     (mm_interconnect_0_key_s1_write),                               //                                           .write
		.KEY_s1_readdata                                  (mm_interconnect_0_key_s1_readdata),                            //                                           .readdata
		.KEY_s1_writedata                                 (mm_interconnect_0_key_s1_writedata),                           //                                           .writedata
		.KEY_s1_chipselect                                (mm_interconnect_0_key_s1_chipselect),                          //                                           .chipselect
		.LCD_DATA_avalon_lcd_slave_address                (mm_interconnect_0_lcd_data_avalon_lcd_slave_address),          //                  LCD_DATA_avalon_lcd_slave.address
		.LCD_DATA_avalon_lcd_slave_write                  (mm_interconnect_0_lcd_data_avalon_lcd_slave_write),            //                                           .write
		.LCD_DATA_avalon_lcd_slave_read                   (mm_interconnect_0_lcd_data_avalon_lcd_slave_read),             //                                           .read
		.LCD_DATA_avalon_lcd_slave_readdata               (mm_interconnect_0_lcd_data_avalon_lcd_slave_readdata),         //                                           .readdata
		.LCD_DATA_avalon_lcd_slave_writedata              (mm_interconnect_0_lcd_data_avalon_lcd_slave_writedata),        //                                           .writedata
		.LCD_DATA_avalon_lcd_slave_waitrequest            (mm_interconnect_0_lcd_data_avalon_lcd_slave_waitrequest),      //                                           .waitrequest
		.LCD_DATA_avalon_lcd_slave_chipselect             (mm_interconnect_0_lcd_data_avalon_lcd_slave_chipselect),       //                                           .chipselect
		.LEDG_s1_address                                  (mm_interconnect_0_ledg_s1_address),                            //                                    LEDG_s1.address
		.LEDG_s1_write                                    (mm_interconnect_0_ledg_s1_write),                              //                                           .write
		.LEDG_s1_readdata                                 (mm_interconnect_0_ledg_s1_readdata),                           //                                           .readdata
		.LEDG_s1_writedata                                (mm_interconnect_0_ledg_s1_writedata),                          //                                           .writedata
		.LEDG_s1_chipselect                               (mm_interconnect_0_ledg_s1_chipselect),                         //                                           .chipselect
		.LEDR_s1_address                                  (mm_interconnect_0_ledr_s1_address),                            //                                    LEDR_s1.address
		.LEDR_s1_write                                    (mm_interconnect_0_ledr_s1_write),                              //                                           .write
		.LEDR_s1_readdata                                 (mm_interconnect_0_ledr_s1_readdata),                           //                                           .readdata
		.LEDR_s1_writedata                                (mm_interconnect_0_ledr_s1_writedata),                          //                                           .writedata
		.LEDR_s1_chipselect                               (mm_interconnect_0_ledr_s1_chipselect),                         //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.on_chip_memory_s1_address                        (mm_interconnect_0_on_chip_memory_s1_address),                  //                          on_chip_memory_s1.address
		.on_chip_memory_s1_write                          (mm_interconnect_0_on_chip_memory_s1_write),                    //                                           .write
		.on_chip_memory_s1_readdata                       (mm_interconnect_0_on_chip_memory_s1_readdata),                 //                                           .readdata
		.on_chip_memory_s1_writedata                      (mm_interconnect_0_on_chip_memory_s1_writedata),                //                                           .writedata
		.on_chip_memory_s1_byteenable                     (mm_interconnect_0_on_chip_memory_s1_byteenable),               //                                           .byteenable
		.on_chip_memory_s1_chipselect                     (mm_interconnect_0_on_chip_memory_s1_chipselect),               //                                           .chipselect
		.on_chip_memory_s1_clken                          (mm_interconnect_0_on_chip_memory_s1_clken),                    //                                           .clken
		.sdram_s1_address                                 (mm_interconnect_0_sdram_s1_address),                           //                                   sdram_s1.address
		.sdram_s1_write                                   (mm_interconnect_0_sdram_s1_write),                             //                                           .write
		.sdram_s1_read                                    (mm_interconnect_0_sdram_s1_read),                              //                                           .read
		.sdram_s1_readdata                                (mm_interconnect_0_sdram_s1_readdata),                          //                                           .readdata
		.sdram_s1_writedata                               (mm_interconnect_0_sdram_s1_writedata),                         //                                           .writedata
		.sdram_s1_byteenable                              (mm_interconnect_0_sdram_s1_byteenable),                        //                                           .byteenable
		.sdram_s1_readdatavalid                           (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                           .readdatavalid
		.sdram_s1_waitrequest                             (mm_interconnect_0_sdram_s1_waitrequest),                       //                                           .waitrequest
		.sdram_s1_chipselect                              (mm_interconnect_0_sdram_s1_chipselect),                        //                                           .chipselect
		.sram_avalon_sram_slave_address                   (mm_interconnect_0_sram_avalon_sram_slave_address),             //                     sram_avalon_sram_slave.address
		.sram_avalon_sram_slave_write                     (mm_interconnect_0_sram_avalon_sram_slave_write),               //                                           .write
		.sram_avalon_sram_slave_read                      (mm_interconnect_0_sram_avalon_sram_slave_read),                //                                           .read
		.sram_avalon_sram_slave_readdata                  (mm_interconnect_0_sram_avalon_sram_slave_readdata),            //                                           .readdata
		.sram_avalon_sram_slave_writedata                 (mm_interconnect_0_sram_avalon_sram_slave_writedata),           //                                           .writedata
		.sram_avalon_sram_slave_byteenable                (mm_interconnect_0_sram_avalon_sram_slave_byteenable),          //                                           .byteenable
		.sram_avalon_sram_slave_readdatavalid             (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),       //                                           .readdatavalid
		.SW_s1_address                                    (mm_interconnect_0_sw_s1_address),                              //                                      SW_s1.address
		.SW_s1_write                                      (mm_interconnect_0_sw_s1_write),                                //                                           .write
		.SW_s1_readdata                                   (mm_interconnect_0_sw_s1_readdata),                             //                                           .readdata
		.SW_s1_writedata                                  (mm_interconnect_0_sw_s1_writedata),                            //                                           .writedata
		.SW_s1_chipselect                                 (mm_interconnect_0_sw_s1_chipselect),                           //                                           .chipselect
		.sysid_qsys_0_control_slave_address               (mm_interconnect_0_sysid_qsys_0_control_slave_address),         //                 sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata              (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),        //                                           .readdata
		.SYSTEM_TIMER_s1_address                          (mm_interconnect_0_system_timer_s1_address),                    //                            SYSTEM_TIMER_s1.address
		.SYSTEM_TIMER_s1_write                            (mm_interconnect_0_system_timer_s1_write),                      //                                           .write
		.SYSTEM_TIMER_s1_readdata                         (mm_interconnect_0_system_timer_s1_readdata),                   //                                           .readdata
		.SYSTEM_TIMER_s1_writedata                        (mm_interconnect_0_system_timer_s1_writedata),                  //                                           .writedata
		.SYSTEM_TIMER_s1_chipselect                       (mm_interconnect_0_system_timer_s1_chipselect)                  //                                           .chipselect
	);

	unsaved_irq_mapper irq_mapper (
		.clk           (clocks_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (clocks_reset_source_reset),                  // reset_in1.reset
		.clk            (clocks_sys_clk_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
